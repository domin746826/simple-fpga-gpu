`ifndef SELECTED_TIMING_VH
`define SELECTED_TIMING_VH

// `include "../timings/800x600.vh"
// `include "../timings/1024x768.vh"
`include "../timings/1440x900.vh"

`endif



