`ifndef VGA_TIMING_1024x768_VH
`define VGA_TIMING_1024x768_VH

// 800x600 @60Hz
`define SMALL_COUNT_TO 4

`define VISIBLE_AREA 1024
`define FRONT_PORCH  24
`define SYNC_PULSE   136
`define BACK_PORCH   160
`define WHOLE_LINE (`VISIBLE_AREA+`FRONT_PORCH+`SYNC_PULSE+`BACK_PORCH)

`define VISIBLE_LINES 768
`define V_FRONT_PORCH 3
`define V_SYNC_PULSE  6
`define V_BACK_PORCH  29
`define WHOLE_FRAME (`VISIBLE_LINES+`V_FRONT_PORCH+`V_SYNC_PULSE+`V_BACK_PORCH)

`define HSYNC_NEGATIVE 1
`define VSYNC_NEGATIVE 1

// 65.000 MHz
`define CLK_DCM_MULTIPLY 13
`define CLK_DCM_DIVIDE   2


// text mode
`define TEXT_COLS 128
`define TEXT_ROWS 48

// graphics mode
`define SIDE_PIXELS_BLACK_GRAPHIC 12
`define BOTTOM_LINES_BLACK_GRAPHIC 18

// text mode
`define SIDE_PIXELS_BLACK_TEXT 0
`define BOTTOM_LINES_BLACK_TEXT 0

`endif
